../SingleCycleProcessor/imem.sv