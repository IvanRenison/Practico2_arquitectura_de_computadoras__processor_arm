/home/ivan/Dropbox/3° 2C Arquitectura del computador/Link to SingleCycleProcessor/execute.sv