../SingleCycleProcessor/fetch.sv