../SingleCycleProcessor/flopr.sv