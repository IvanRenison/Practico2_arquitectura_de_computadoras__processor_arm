../SingleCycleProcessor/signext.sv