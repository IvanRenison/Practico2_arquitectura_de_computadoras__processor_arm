../SingleCycleProcessor/regfile.sv