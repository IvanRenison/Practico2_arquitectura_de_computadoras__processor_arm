../SingleCycleProcessor/adder.sv