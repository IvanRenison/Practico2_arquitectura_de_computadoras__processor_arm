../SingleCycleProcessor/execute.sv