../SingleCycleProcessor/alu.sv