../SingleCycleProcessor/maindec.sv